interface spi_interface;
    logic sck_o; //serial clk
    logic miso_i; //master in
    logic mosi_o; //master out
endinterface e spi_interface