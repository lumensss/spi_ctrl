class className;
    function new();
        
    endfunction //new()
endclass //className