//  Class: cdn_cdrlftest 
//
class cdn_cdrlftest extends uvm_agent;
    //  Group: Variables


    //  Group: Constraints


    //  Group: Functions

    //  Constructor: new
    function new(string name = "cdn_cdrlftest ");
    endfunction: new
    

endclass: cdn_cdrlftest 
